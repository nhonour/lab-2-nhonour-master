module task4(input logic CLOCK_50, input logic KEY[3:0], // KEY[3] is async active-low reset
             output logic [9:0] VGA_R, output logic [9:0] VGA_G, output logic [9:0] VGA_B,
             output logic VGA_HS, output logic VGA_VS,
             output logic VGA_BLANK, output logic VGA_SYNC, output logic VGA_CLK);
  
    // instantiate and connect the VGA adapter and your module

endmodule

