module filledcircle(input logic clk, input logic rstn, input logic [2:0] colour,
                    input logic [7:0] centre_x, input logic [6:0] centre_y, input logic [7:0] radius,
                    input logic start, output logic done,
                    output logic [7:0] vga_x, output logic [6:0] vga_y,
                    output logic [2:0] vga_colour, output logic vga_plot);
     // draw the filled circle
endmodule

